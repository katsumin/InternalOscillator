// megafunction wizard: %MAX II/MAX V oscillator%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTUFM_OSC 

// ============================================================
// File Name: osc.v
// Megafunction Name(s):
// 			ALTUFM_OSC
//
// Simulation Library Files(s):
// 			maxv
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// ************************************************************

//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.

module osc (
	oscena,
	osc)/* synthesis synthesis_clearbox = 1 */;

	input	  oscena;
	output	  osc;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX V"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altufm_osc"
// Retrieval info: CONSTANT: OSC_FREQUENCY NUMERIC "188679"
// Retrieval info: USED_PORT: osc 0 0 0 0 OUTPUT NODEFVAL "osc"
// Retrieval info: CONNECT: osc 0 0 0 0 @osc 0 0 0 0
// Retrieval info: USED_PORT: oscena 0 0 0 0 INPUT NODEFVAL "oscena"
// Retrieval info: CONNECT: @oscena 0 0 0 0 oscena 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL osc.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL osc.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL osc.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL osc_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL osc_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL osc.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL osc.cmp TRUE TRUE
// Retrieval info: LIB_FILE: maxv
